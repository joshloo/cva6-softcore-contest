component osc0 is
    port(
        en_i: in std_logic;
        clk_sel_i: in std_logic;
        clk_out_o: out std_logic
    );
end component;

__: osc0 port map(
    en_i=>,
    clk_sel_i=>,
    clk_out_o=>
);
